module test;
endmodule